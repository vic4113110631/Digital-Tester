// Architectire.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module Architectire (
		input  wire        clk_clk,                                       //                           clk.clk
		output wire        clockbridge_out_clk,                           //               clockbridge_out.clk
		output wire        controlsignal_export,                          //                 controlsignal.export
		input  wire        dcfifo_csr_address,                            //                    dcfifo_csr.address
		input  wire        dcfifo_csr_read,                               //                              .read
		input  wire        dcfifo_csr_write,                              //                              .write
		output wire [31:0] dcfifo_csr_readdata,                           //                              .readdata
		input  wire [31:0] dcfifo_csr_writedata,                          //                              .writedata
		output wire [31:0] dcfifo_out_data,                               //                    dcfifo_out.data
		output wire        dcfifo_out_valid,                              //                              .valid
		input  wire        dcfifo_out_ready,                              //                              .ready
		output wire        dcfifo_out_startofpacket,                      //                              .startofpacket
		output wire        dcfifo_out_endofpacket,                        //                              .endofpacket
		output wire        pciexpress_clocks_sim_clk250_export,           //         pciexpress_clocks_sim.clk250_export
		output wire        pciexpress_clocks_sim_clk500_export,           //                              .clk500_export
		output wire        pciexpress_clocks_sim_clk125_export,           //                              .clk125_export
		input  wire        pciexpress_pipe_ext_pipe_mode,                 //           pciexpress_pipe_ext.pipe_mode
		input  wire        pciexpress_pipe_ext_phystatus_ext,             //                              .phystatus_ext
		output wire        pciexpress_pipe_ext_rate_ext,                  //                              .rate_ext
		output wire [1:0]  pciexpress_pipe_ext_powerdown_ext,             //                              .powerdown_ext
		output wire        pciexpress_pipe_ext_txdetectrx_ext,            //                              .txdetectrx_ext
		input  wire        pciexpress_pipe_ext_rxelecidle0_ext,           //                              .rxelecidle0_ext
		input  wire [7:0]  pciexpress_pipe_ext_rxdata0_ext,               //                              .rxdata0_ext
		input  wire [2:0]  pciexpress_pipe_ext_rxstatus0_ext,             //                              .rxstatus0_ext
		input  wire        pciexpress_pipe_ext_rxvalid0_ext,              //                              .rxvalid0_ext
		input  wire        pciexpress_pipe_ext_rxdatak0_ext,              //                              .rxdatak0_ext
		output wire [7:0]  pciexpress_pipe_ext_txdata0_ext,               //                              .txdata0_ext
		output wire        pciexpress_pipe_ext_txdatak0_ext,              //                              .txdatak0_ext
		output wire        pciexpress_pipe_ext_rxpolarity0_ext,           //                              .rxpolarity0_ext
		output wire        pciexpress_pipe_ext_txcompl0_ext,              //                              .txcompl0_ext
		output wire        pciexpress_pipe_ext_txelecidle0_ext,           //                              .txelecidle0_ext
		input  wire        pciexpress_powerdown_pll_powerdown,            //          pciexpress_powerdown.pll_powerdown
		input  wire        pciexpress_powerdown_gxb_powerdown,            //                              .gxb_powerdown
		input  wire        pciexpress_reconfig_busy_busy_altgxb_reconfig, //      pciexpress_reconfig_busy.busy_altgxb_reconfig
		output wire [4:0]  pciexpress_reconfig_fromgxb_0_data,            // pciexpress_reconfig_fromgxb_0.data
		input  wire [3:0]  pciexpress_reconfig_togxb_data,                //     pciexpress_reconfig_togxb.data
		input  wire        pciexpress_refclk_export,                      //             pciexpress_refclk.export
		input  wire        pciexpress_rstn_export,                        //               pciexpress_rstn.export
		input  wire        pciexpress_rx_in_rx_datain_0,                  //              pciexpress_rx_in.rx_datain_0
		input  wire [39:0] pciexpress_test_in_test_in,                    //            pciexpress_test_in.test_in
		output wire        pciexpress_tx_out_tx_dataout_0,                //             pciexpress_tx_out.tx_dataout_0
		input  wire        reset_reset_n,                                 //                         reset.reset_n
		input  wire [10:0] response_export                                //                      response.export
	);

	wire         pll_c0_clk;                                     // PLL:c0 -> [PCIExpress:cal_blk_clk_clk, PCIExpress:reconfig_gxbclk_clk]
	wire         pciexpress_pcie_core_clk_clk;                   // PCIExpress:pcie_core_clk_clk -> [ControlSignal:clk, DCFIFO:in_clk, FIFO_Memory:wrclock, PCIExpress:fixedclk_clk, Response:clk, SGDMA:clk, avalon_st_adapter:in_clk_0_clk, irq_mapper:clk, mm_interconnect_0:PCIExpress_pcie_core_clk_clk, mm_interconnect_1:PCIExpress_pcie_core_clk_clk, mm_interconnect_2:PCIExpress_pcie_core_clk_clk, rst_controller:clk, rst_controller_001:clk]
	wire         pciexpress_bar1_0_waitrequest;                  // mm_interconnect_0:PCIExpress_bar1_0_waitrequest -> PCIExpress:bar1_0_waitrequest
	wire  [63:0] pciexpress_bar1_0_readdata;                     // mm_interconnect_0:PCIExpress_bar1_0_readdata -> PCIExpress:bar1_0_readdata
	wire  [31:0] pciexpress_bar1_0_address;                      // PCIExpress:bar1_0_address -> mm_interconnect_0:PCIExpress_bar1_0_address
	wire         pciexpress_bar1_0_read;                         // PCIExpress:bar1_0_read -> mm_interconnect_0:PCIExpress_bar1_0_read
	wire   [7:0] pciexpress_bar1_0_byteenable;                   // PCIExpress:bar1_0_byteenable -> mm_interconnect_0:PCIExpress_bar1_0_byteenable
	wire         pciexpress_bar1_0_readdatavalid;                // mm_interconnect_0:PCIExpress_bar1_0_readdatavalid -> PCIExpress:bar1_0_readdatavalid
	wire         pciexpress_bar1_0_write;                        // PCIExpress:bar1_0_write -> mm_interconnect_0:PCIExpress_bar1_0_write
	wire  [63:0] pciexpress_bar1_0_writedata;                    // PCIExpress:bar1_0_writedata -> mm_interconnect_0:PCIExpress_bar1_0_writedata
	wire   [6:0] pciexpress_bar1_0_burstcount;                   // PCIExpress:bar1_0_burstcount -> mm_interconnect_0:PCIExpress_bar1_0_burstcount
	wire         sgdma_m_write_waitrequest;                      // mm_interconnect_0:SGDMA_m_write_waitrequest -> SGDMA:m_write_waitrequest
	wire  [31:0] sgdma_m_write_address;                          // SGDMA:m_write_address -> mm_interconnect_0:SGDMA_m_write_address
	wire   [3:0] sgdma_m_write_byteenable;                       // SGDMA:m_write_byteenable -> mm_interconnect_0:SGDMA_m_write_byteenable
	wire         sgdma_m_write_write;                            // SGDMA:m_write_write -> mm_interconnect_0:SGDMA_m_write_write
	wire  [31:0] sgdma_m_write_writedata;                        // SGDMA:m_write_writedata -> mm_interconnect_0:SGDMA_m_write_writedata
	wire         mm_interconnect_0_fifo_memory_in_waitrequest;   // FIFO_Memory:avalonmm_write_slave_waitrequest -> mm_interconnect_0:FIFO_Memory_in_waitrequest
	wire   [0:0] mm_interconnect_0_fifo_memory_in_address;       // mm_interconnect_0:FIFO_Memory_in_address -> FIFO_Memory:avalonmm_write_slave_address
	wire         mm_interconnect_0_fifo_memory_in_write;         // mm_interconnect_0:FIFO_Memory_in_write -> FIFO_Memory:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_memory_in_writedata;     // mm_interconnect_0:FIFO_Memory_in_writedata -> FIFO_Memory:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_response_s1_readdata;         // Response:readdata -> mm_interconnect_0:Response_s1_readdata
	wire   [1:0] mm_interconnect_0_response_s1_address;          // mm_interconnect_0:Response_s1_address -> Response:address
	wire         mm_interconnect_0_controlsignal_s1_chipselect;  // mm_interconnect_0:ControlSignal_s1_chipselect -> ControlSignal:chipselect
	wire  [31:0] mm_interconnect_0_controlsignal_s1_readdata;    // ControlSignal:readdata -> mm_interconnect_0:ControlSignal_s1_readdata
	wire   [1:0] mm_interconnect_0_controlsignal_s1_address;     // mm_interconnect_0:ControlSignal_s1_address -> ControlSignal:address
	wire         mm_interconnect_0_controlsignal_s1_write;       // mm_interconnect_0:ControlSignal_s1_write -> ControlSignal:write_n
	wire  [31:0] mm_interconnect_0_controlsignal_s1_writedata;   // mm_interconnect_0:ControlSignal_s1_writedata -> ControlSignal:writedata
	wire         pciexpress_bar2_waitrequest;                    // mm_interconnect_1:PCIExpress_bar2_waitrequest -> PCIExpress:bar2_waitrequest
	wire  [63:0] pciexpress_bar2_readdata;                       // mm_interconnect_1:PCIExpress_bar2_readdata -> PCIExpress:bar2_readdata
	wire  [31:0] pciexpress_bar2_address;                        // PCIExpress:bar2_address -> mm_interconnect_1:PCIExpress_bar2_address
	wire         pciexpress_bar2_read;                           // PCIExpress:bar2_read -> mm_interconnect_1:PCIExpress_bar2_read
	wire   [7:0] pciexpress_bar2_byteenable;                     // PCIExpress:bar2_byteenable -> mm_interconnect_1:PCIExpress_bar2_byteenable
	wire         pciexpress_bar2_readdatavalid;                  // mm_interconnect_1:PCIExpress_bar2_readdatavalid -> PCIExpress:bar2_readdatavalid
	wire         pciexpress_bar2_write;                          // PCIExpress:bar2_write -> mm_interconnect_1:PCIExpress_bar2_write
	wire  [63:0] pciexpress_bar2_writedata;                      // PCIExpress:bar2_writedata -> mm_interconnect_1:PCIExpress_bar2_writedata
	wire   [6:0] pciexpress_bar2_burstcount;                     // PCIExpress:bar2_burstcount -> mm_interconnect_1:PCIExpress_bar2_burstcount
	wire         mm_interconnect_1_pciexpress_cra_chipselect;    // mm_interconnect_1:PCIExpress_cra_chipselect -> PCIExpress:cra_chipselect
	wire  [31:0] mm_interconnect_1_pciexpress_cra_readdata;      // PCIExpress:cra_readdata -> mm_interconnect_1:PCIExpress_cra_readdata
	wire         mm_interconnect_1_pciexpress_cra_waitrequest;   // PCIExpress:cra_waitrequest -> mm_interconnect_1:PCIExpress_cra_waitrequest
	wire  [11:0] mm_interconnect_1_pciexpress_cra_address;       // mm_interconnect_1:PCIExpress_cra_address -> PCIExpress:cra_address
	wire         mm_interconnect_1_pciexpress_cra_read;          // mm_interconnect_1:PCIExpress_cra_read -> PCIExpress:cra_read
	wire   [3:0] mm_interconnect_1_pciexpress_cra_byteenable;    // mm_interconnect_1:PCIExpress_cra_byteenable -> PCIExpress:cra_byteenable
	wire         mm_interconnect_1_pciexpress_cra_write;         // mm_interconnect_1:PCIExpress_cra_write -> PCIExpress:cra_write
	wire  [31:0] mm_interconnect_1_pciexpress_cra_writedata;     // mm_interconnect_1:PCIExpress_cra_writedata -> PCIExpress:cra_writedata
	wire         mm_interconnect_1_sgdma_csr_chipselect;         // mm_interconnect_1:SGDMA_csr_chipselect -> SGDMA:csr_chipselect
	wire  [31:0] mm_interconnect_1_sgdma_csr_readdata;           // SGDMA:csr_readdata -> mm_interconnect_1:SGDMA_csr_readdata
	wire   [3:0] mm_interconnect_1_sgdma_csr_address;            // mm_interconnect_1:SGDMA_csr_address -> SGDMA:csr_address
	wire         mm_interconnect_1_sgdma_csr_read;               // mm_interconnect_1:SGDMA_csr_read -> SGDMA:csr_read
	wire         mm_interconnect_1_sgdma_csr_write;              // mm_interconnect_1:SGDMA_csr_write -> SGDMA:csr_write
	wire  [31:0] mm_interconnect_1_sgdma_csr_writedata;          // mm_interconnect_1:SGDMA_csr_writedata -> SGDMA:csr_writedata
	wire  [31:0] sgdma_descriptor_read_readdata;                 // mm_interconnect_2:SGDMA_descriptor_read_readdata -> SGDMA:descriptor_read_readdata
	wire         sgdma_descriptor_read_waitrequest;              // mm_interconnect_2:SGDMA_descriptor_read_waitrequest -> SGDMA:descriptor_read_waitrequest
	wire  [31:0] sgdma_descriptor_read_address;                  // SGDMA:descriptor_read_address -> mm_interconnect_2:SGDMA_descriptor_read_address
	wire         sgdma_descriptor_read_read;                     // SGDMA:descriptor_read_read -> mm_interconnect_2:SGDMA_descriptor_read_read
	wire         sgdma_descriptor_read_readdatavalid;            // mm_interconnect_2:SGDMA_descriptor_read_readdatavalid -> SGDMA:descriptor_read_readdatavalid
	wire         sgdma_descriptor_write_waitrequest;             // mm_interconnect_2:SGDMA_descriptor_write_waitrequest -> SGDMA:descriptor_write_waitrequest
	wire  [31:0] sgdma_descriptor_write_address;                 // SGDMA:descriptor_write_address -> mm_interconnect_2:SGDMA_descriptor_write_address
	wire         sgdma_descriptor_write_write;                   // SGDMA:descriptor_write_write -> mm_interconnect_2:SGDMA_descriptor_write_write
	wire  [31:0] sgdma_descriptor_write_writedata;               // SGDMA:descriptor_write_writedata -> mm_interconnect_2:SGDMA_descriptor_write_writedata
	wire  [31:0] sgdma_m_read_readdata;                          // mm_interconnect_2:SGDMA_m_read_readdata -> SGDMA:m_read_readdata
	wire         sgdma_m_read_waitrequest;                       // mm_interconnect_2:SGDMA_m_read_waitrequest -> SGDMA:m_read_waitrequest
	wire  [31:0] sgdma_m_read_address;                           // SGDMA:m_read_address -> mm_interconnect_2:SGDMA_m_read_address
	wire         sgdma_m_read_read;                              // SGDMA:m_read_read -> mm_interconnect_2:SGDMA_m_read_read
	wire         sgdma_m_read_readdatavalid;                     // mm_interconnect_2:SGDMA_m_read_readdatavalid -> SGDMA:m_read_readdatavalid
	wire         mm_interconnect_2_pciexpress_txs_chipselect;    // mm_interconnect_2:PCIExpress_txs_chipselect -> PCIExpress:txs_chipselect
	wire  [63:0] mm_interconnect_2_pciexpress_txs_readdata;      // PCIExpress:txs_readdata -> mm_interconnect_2:PCIExpress_txs_readdata
	wire         mm_interconnect_2_pciexpress_txs_waitrequest;   // PCIExpress:txs_waitrequest -> mm_interconnect_2:PCIExpress_txs_waitrequest
	wire  [30:0] mm_interconnect_2_pciexpress_txs_address;       // mm_interconnect_2:PCIExpress_txs_address -> PCIExpress:txs_address
	wire         mm_interconnect_2_pciexpress_txs_read;          // mm_interconnect_2:PCIExpress_txs_read -> PCIExpress:txs_read
	wire   [7:0] mm_interconnect_2_pciexpress_txs_byteenable;    // mm_interconnect_2:PCIExpress_txs_byteenable -> PCIExpress:txs_byteenable
	wire         mm_interconnect_2_pciexpress_txs_readdatavalid; // PCIExpress:txs_readdatavalid -> mm_interconnect_2:PCIExpress_txs_readdatavalid
	wire         mm_interconnect_2_pciexpress_txs_write;         // mm_interconnect_2:PCIExpress_txs_write -> PCIExpress:txs_write
	wire  [63:0] mm_interconnect_2_pciexpress_txs_writedata;     // mm_interconnect_2:PCIExpress_txs_writedata -> PCIExpress:txs_writedata
	wire   [6:0] mm_interconnect_2_pciexpress_txs_burstcount;    // mm_interconnect_2:PCIExpress_txs_burstcount -> PCIExpress:txs_burstcount
	wire         irq_mapper_receiver0_irq;                       // SGDMA:csr_irq -> irq_mapper:receiver0_irq
	wire  [15:0] pciexpress_rxm_irq_irq;                         // irq_mapper:sender_irq -> PCIExpress:rxm_irq_irq
	wire         fifo_memory_out_valid;                          // FIFO_Memory:avalonst_source_valid -> avalon_st_adapter:in_0_valid
	wire  [31:0] fifo_memory_out_data;                           // FIFO_Memory:avalonst_source_data -> avalon_st_adapter:in_0_data
	wire         fifo_memory_out_ready;                          // avalon_st_adapter:in_0_ready -> FIFO_Memory:avalonst_source_ready
	wire   [7:0] fifo_memory_out_channel;                        // FIFO_Memory:avalonst_source_channel -> avalon_st_adapter:in_0_channel
	wire         fifo_memory_out_startofpacket;                  // FIFO_Memory:avalonst_source_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire   [7:0] fifo_memory_out_error;                          // FIFO_Memory:avalonst_source_error -> avalon_st_adapter:in_0_error
	wire         fifo_memory_out_endofpacket;                    // FIFO_Memory:avalonst_source_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                  // avalon_st_adapter:out_0_valid -> DCFIFO:in_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                   // avalon_st_adapter:out_0_data -> DCFIFO:in_data
	wire         avalon_st_adapter_out_0_ready;                  // DCFIFO:in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;          // avalon_st_adapter:out_0_startofpacket -> DCFIFO:in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;            // avalon_st_adapter:out_0_endofpacket -> DCFIFO:in_endofpacket
	wire         rst_controller_reset_out_reset;                 // rst_controller:reset_out -> [ControlSignal:reset_n, FIFO_Memory:reset_n, Response:reset_n, SGDMA:system_reset_n, avalon_st_adapter:in_rst_0_reset, mm_interconnect_0:SGDMA_reset_reset_bridge_in_reset_reset, mm_interconnect_1:SGDMA_reset_reset_bridge_in_reset_reset, mm_interconnect_2:SGDMA_reset_reset_bridge_in_reset_reset]
	wire         pciexpress_pcie_core_reset_reset;               // PCIExpress:pcie_core_reset_reset_n -> [rst_controller:reset_in1, rst_controller_001:reset_in0, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;             // rst_controller_001:reset_out -> [DCFIFO:in_reset_n, irq_mapper:reset, mm_interconnect_0:PCIExpress_bar1_0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:PCIExpress_bar2_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:PCIExpress_txs_translator_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;             // rst_controller_002:reset_out -> DCFIFO:out_reset_n
	wire         rst_controller_003_reset_out_reset;             // rst_controller_003:reset_out -> PLL:reset

	Architectire_ControlSignal controlsignal (
		.clk        (pciexpress_pcie_core_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_controlsignal_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_controlsignal_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_controlsignal_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_controlsignal_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_controlsignal_s1_readdata),   //                    .readdata
		.out_port   (controlsignal_export)                           // external_connection.export
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (1),
		.BITS_PER_SYMBOL    (32),
		.FIFO_DEPTH         (65536),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (1),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (1),
		.WR_SYNC_DEPTH      (32),
		.RD_SYNC_DEPTH      (32)
	) dcfifo (
		.in_clk            (pciexpress_pcie_core_clk_clk),          //        in_clk.clk
		.in_reset_n        (~rst_controller_001_reset_out_reset),   //  in_clk_reset.reset_n
		.out_clk           (clockbridge_out_clk),                   //       out_clk.clk
		.out_reset_n       (~rst_controller_002_reset_out_reset),   // out_clk_reset.reset_n
		.out_csr_address   (dcfifo_csr_address),                    //       out_csr.address
		.out_csr_read      (dcfifo_csr_read),                       //              .read
		.out_csr_write     (dcfifo_csr_write),                      //              .write
		.out_csr_readdata  (dcfifo_csr_readdata),                   //              .readdata
		.out_csr_writedata (dcfifo_csr_writedata),                  //              .writedata
		.in_data           (avalon_st_adapter_out_0_data),          //            in.data
		.in_valid          (avalon_st_adapter_out_0_valid),         //              .valid
		.in_ready          (avalon_st_adapter_out_0_ready),         //              .ready
		.in_startofpacket  (avalon_st_adapter_out_0_startofpacket), //              .startofpacket
		.in_endofpacket    (avalon_st_adapter_out_0_endofpacket),   //              .endofpacket
		.out_data          (dcfifo_out_data),                       //           out.data
		.out_valid         (dcfifo_out_valid),                      //              .valid
		.out_ready         (dcfifo_out_ready),                      //              .ready
		.out_startofpacket (dcfifo_out_startofpacket),              //              .startofpacket
		.out_endofpacket   (dcfifo_out_endofpacket),                //              .endofpacket
		.in_csr_address    (1'b0),                                  //   (terminated)
		.in_csr_read       (1'b0),                                  //   (terminated)
		.in_csr_write      (1'b0),                                  //   (terminated)
		.in_csr_readdata   (),                                      //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000)   //   (terminated)
	);

	Architectire_FIFO_Memory fifo_memory (
		.wrclock                          (pciexpress_pcie_core_clk_clk),                 //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),              // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_memory_in_writedata),   //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_memory_in_write),       //         .write
		.avalonmm_write_slave_address     (mm_interconnect_0_fifo_memory_in_address),     //         .address
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_memory_in_waitrequest), //         .waitrequest
		.avalonst_source_valid            (fifo_memory_out_valid),                        //      out.valid
		.avalonst_source_data             (fifo_memory_out_data),                         //         .data
		.avalonst_source_channel          (fifo_memory_out_channel),                      //         .channel
		.avalonst_source_error            (fifo_memory_out_error),                        //         .error
		.avalonst_source_startofpacket    (fifo_memory_out_startofpacket),                //         .startofpacket
		.avalonst_source_endofpacket      (fifo_memory_out_endofpacket),                  //         .endofpacket
		.avalonst_source_ready            (fifo_memory_out_ready)                         //         .ready
	);

	Architectire_PCIExpress #(
		.p_pcie_hip_type                     ("2"),
		.lane_mask                           (8'b11111110),
		.max_link_width                      (1),
		.millisecond_cycle_count             ("125000"),
		.enable_gen2_core                    ("false"),
		.gen2_lane_rate_mode                 ("false"),
		.no_soft_reset                       ("false"),
		.core_clk_divider                    (2),
		.enable_ch0_pclk_out                 ("true"),
		.core_clk_source                     ("pclk"),
		.CB_P2A_AVALON_ADDR_B0               (0),
		.bar0_size_mask                      (6),
		.bar0_io_space                       ("false"),
		.bar0_64bit_mem_space                ("true"),
		.bar0_prefetchable                   ("true"),
		.CB_P2A_AVALON_ADDR_B1               (0),
		.bar1_size_mask                      (0),
		.bar1_io_space                       ("false"),
		.bar1_64bit_mem_space                ("true"),
		.bar1_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B2               (0),
		.bar2_size_mask                      (15),
		.bar2_io_space                       ("false"),
		.bar2_64bit_mem_space                ("false"),
		.bar2_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B3               (0),
		.bar3_size_mask                      (0),
		.bar3_io_space                       ("false"),
		.bar3_64bit_mem_space                ("false"),
		.bar3_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B4               (0),
		.bar4_size_mask                      (0),
		.bar4_io_space                       ("false"),
		.bar4_64bit_mem_space                ("false"),
		.bar4_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B5               (0),
		.bar5_size_mask                      (0),
		.bar5_io_space                       ("false"),
		.bar5_64bit_mem_space                ("false"),
		.bar5_prefetchable                   ("false"),
		.vendor_id                           (4466),
		.device_id                           (57345),
		.revision_id                         (1),
		.class_code                          (0),
		.subsystem_vendor_id                 (4466),
		.subsystem_device_id                 (4),
		.port_link_number                    (1),
		.msi_function_count                  (0),
		.enable_msi_64bit_addressing         ("true"),
		.enable_function_msix_support        ("false"),
		.eie_before_nfts_count               (4),
		.enable_completion_timeout_disable   ("false"),
		.completion_timeout                  ("NONE"),
		.enable_adapter_half_rate_mode       ("false"),
		.msix_pba_bir                        (0),
		.msix_pba_offset                     (0),
		.msix_table_bir                      (0),
		.msix_table_offset                   (0),
		.msix_table_size                     (0),
		.use_crc_forwarding                  ("false"),
		.surprise_down_error_support         ("false"),
		.dll_active_report_support           ("false"),
		.bar_io_window_size                  ("32BIT"),
		.bar_prefetchable                    (32),
		.hot_plug_support                    (7'b0000000),
		.no_command_completed                ("true"),
		.slot_power_limit                    (0),
		.slot_power_scale                    (0),
		.slot_number                         (0),
		.enable_slot_register                ("false"),
		.advanced_errors                     ("false"),
		.enable_ecrc_check                   ("false"),
		.enable_ecrc_gen                     ("false"),
		.max_payload_size                    (1),
		.retry_buffer_last_active_address    (255),
		.credit_buffer_allocation_aux        ("ABSOLUTE"),
		.vc0_rx_flow_ctrl_posted_header      (28),
		.vc0_rx_flow_ctrl_posted_data        (198),
		.vc0_rx_flow_ctrl_nonposted_header   (30),
		.vc0_rx_flow_ctrl_nonposted_data     (0),
		.vc0_rx_flow_ctrl_compl_header       (48),
		.vc0_rx_flow_ctrl_compl_data         (256),
		.RX_BUF                              (9),
		.RH_NUM                              (7),
		.G_TAG_NUM0                          (32),
		.endpoint_l0_latency                 (0),
		.endpoint_l1_latency                 (0),
		.enable_l1_aspm                      ("false"),
		.l01_entry_latency                   (31),
		.diffclock_nfts_count                (255),
		.sameclock_nfts_count                (255),
		.l1_exit_latency_sameclock           (7),
		.l1_exit_latency_diffclock           (7),
		.l0_exit_latency_sameclock           (7),
		.l0_exit_latency_diffclock           (7),
		.gen2_diffclock_nfts_count           (255),
		.gen2_sameclock_nfts_count           (255),
		.CG_COMMON_CLOCK_MODE                (1),
		.CB_PCIE_MODE                        (0),
		.AST_LITE                            (0),
		.CB_PCIE_RX_LITE                     (0),
		.CG_RXM_IRQ_NUM                      (16),
		.CG_AVALON_S_ADDR_WIDTH              (20),
		.bypass_tl                           ("false"),
		.CG_IMPL_CRA_AV_SLAVE_PORT           (1),
		.CG_NO_CPL_REORDERING                (0),
		.CG_ENABLE_A2P_INTERRUPT             (0),
		.p_user_msi_enable                   (0),
		.CG_IRQ_BIT_ENA                      (65535),
		.CB_A2P_ADDR_MAP_IS_FIXED            (1),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES         (1),
		.CB_A2P_ADDR_MAP_PASS_THRU_BITS      (31),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_LOW  (32'b00000000000000000000000000000000),
		.RXM_DATA_WIDTH                      (64),
		.RXM_BEN_WIDTH                       (8),
		.TL_SELECTION                        (1),
		.pcie_mode                           ("SHARED_MODE"),
		.single_rx_detect                    (1),
		.enable_coreclk_out_half_rate        ("false"),
		.low_priority_vc                     (0),
		.link_width                          (1),
		.cyclone4                            (1)
	) pciexpress (
		.pcie_core_clk_clk                  (pciexpress_pcie_core_clk_clk),                   //      pcie_core_clk.clk
		.pcie_core_reset_reset_n            (pciexpress_pcie_core_reset_reset),               //    pcie_core_reset.reset_n
		.cal_blk_clk_clk                    (pll_c0_clk),                                     //        cal_blk_clk.clk
		.txs_address                        (mm_interconnect_2_pciexpress_txs_address),       //                txs.address
		.txs_chipselect                     (mm_interconnect_2_pciexpress_txs_chipselect),    //                   .chipselect
		.txs_byteenable                     (mm_interconnect_2_pciexpress_txs_byteenable),    //                   .byteenable
		.txs_readdata                       (mm_interconnect_2_pciexpress_txs_readdata),      //                   .readdata
		.txs_writedata                      (mm_interconnect_2_pciexpress_txs_writedata),     //                   .writedata
		.txs_read                           (mm_interconnect_2_pciexpress_txs_read),          //                   .read
		.txs_write                          (mm_interconnect_2_pciexpress_txs_write),         //                   .write
		.txs_burstcount                     (mm_interconnect_2_pciexpress_txs_burstcount),    //                   .burstcount
		.txs_readdatavalid                  (mm_interconnect_2_pciexpress_txs_readdatavalid), //                   .readdatavalid
		.txs_waitrequest                    (mm_interconnect_2_pciexpress_txs_waitrequest),   //                   .waitrequest
		.refclk_export                      (pciexpress_refclk_export),                       //             refclk.export
		.test_in_test_in                    (pciexpress_test_in_test_in),                     //            test_in.test_in
		.pcie_rstn_export                   (pciexpress_rstn_export),                         //          pcie_rstn.export
		.clocks_sim_clk250_export           (pciexpress_clocks_sim_clk250_export),            //         clocks_sim.clk250_export
		.clocks_sim_clk500_export           (pciexpress_clocks_sim_clk500_export),            //                   .clk500_export
		.clocks_sim_clk125_export           (pciexpress_clocks_sim_clk125_export),            //                   .clk125_export
		.reconfig_busy_busy_altgxb_reconfig (pciexpress_reconfig_busy_busy_altgxb_reconfig),  //      reconfig_busy.busy_altgxb_reconfig
		.pipe_ext_pipe_mode                 (pciexpress_pipe_ext_pipe_mode),                  //           pipe_ext.pipe_mode
		.pipe_ext_phystatus_ext             (pciexpress_pipe_ext_phystatus_ext),              //                   .phystatus_ext
		.pipe_ext_rate_ext                  (pciexpress_pipe_ext_rate_ext),                   //                   .rate_ext
		.pipe_ext_powerdown_ext             (pciexpress_pipe_ext_powerdown_ext),              //                   .powerdown_ext
		.pipe_ext_txdetectrx_ext            (pciexpress_pipe_ext_txdetectrx_ext),             //                   .txdetectrx_ext
		.pipe_ext_rxelecidle0_ext           (pciexpress_pipe_ext_rxelecidle0_ext),            //                   .rxelecidle0_ext
		.pipe_ext_rxdata0_ext               (pciexpress_pipe_ext_rxdata0_ext),                //                   .rxdata0_ext
		.pipe_ext_rxstatus0_ext             (pciexpress_pipe_ext_rxstatus0_ext),              //                   .rxstatus0_ext
		.pipe_ext_rxvalid0_ext              (pciexpress_pipe_ext_rxvalid0_ext),               //                   .rxvalid0_ext
		.pipe_ext_rxdatak0_ext              (pciexpress_pipe_ext_rxdatak0_ext),               //                   .rxdatak0_ext
		.pipe_ext_txdata0_ext               (pciexpress_pipe_ext_txdata0_ext),                //                   .txdata0_ext
		.pipe_ext_txdatak0_ext              (pciexpress_pipe_ext_txdatak0_ext),               //                   .txdatak0_ext
		.pipe_ext_rxpolarity0_ext           (pciexpress_pipe_ext_rxpolarity0_ext),            //                   .rxpolarity0_ext
		.pipe_ext_txcompl0_ext              (pciexpress_pipe_ext_txcompl0_ext),               //                   .txcompl0_ext
		.pipe_ext_txelecidle0_ext           (pciexpress_pipe_ext_txelecidle0_ext),            //                   .txelecidle0_ext
		.powerdown_pll_powerdown            (pciexpress_powerdown_pll_powerdown),             //          powerdown.pll_powerdown
		.powerdown_gxb_powerdown            (pciexpress_powerdown_gxb_powerdown),             //                   .gxb_powerdown
		.bar1_0_address                     (pciexpress_bar1_0_address),                      //             bar1_0.address
		.bar1_0_read                        (pciexpress_bar1_0_read),                         //                   .read
		.bar1_0_waitrequest                 (pciexpress_bar1_0_waitrequest),                  //                   .waitrequest
		.bar1_0_write                       (pciexpress_bar1_0_write),                        //                   .write
		.bar1_0_readdatavalid               (pciexpress_bar1_0_readdatavalid),                //                   .readdatavalid
		.bar1_0_readdata                    (pciexpress_bar1_0_readdata),                     //                   .readdata
		.bar1_0_writedata                   (pciexpress_bar1_0_writedata),                    //                   .writedata
		.bar1_0_burstcount                  (pciexpress_bar1_0_burstcount),                   //                   .burstcount
		.bar1_0_byteenable                  (pciexpress_bar1_0_byteenable),                   //                   .byteenable
		.bar2_address                       (pciexpress_bar2_address),                        //               bar2.address
		.bar2_read                          (pciexpress_bar2_read),                           //                   .read
		.bar2_waitrequest                   (pciexpress_bar2_waitrequest),                    //                   .waitrequest
		.bar2_write                         (pciexpress_bar2_write),                          //                   .write
		.bar2_readdatavalid                 (pciexpress_bar2_readdatavalid),                  //                   .readdatavalid
		.bar2_readdata                      (pciexpress_bar2_readdata),                       //                   .readdata
		.bar2_writedata                     (pciexpress_bar2_writedata),                      //                   .writedata
		.bar2_burstcount                    (pciexpress_bar2_burstcount),                     //                   .burstcount
		.bar2_byteenable                    (pciexpress_bar2_byteenable),                     //                   .byteenable
		.cra_chipselect                     (mm_interconnect_1_pciexpress_cra_chipselect),    //                cra.chipselect
		.cra_address                        (mm_interconnect_1_pciexpress_cra_address),       //                   .address
		.cra_byteenable                     (mm_interconnect_1_pciexpress_cra_byteenable),    //                   .byteenable
		.cra_read                           (mm_interconnect_1_pciexpress_cra_read),          //                   .read
		.cra_readdata                       (mm_interconnect_1_pciexpress_cra_readdata),      //                   .readdata
		.cra_write                          (mm_interconnect_1_pciexpress_cra_write),         //                   .write
		.cra_writedata                      (mm_interconnect_1_pciexpress_cra_writedata),     //                   .writedata
		.cra_waitrequest                    (mm_interconnect_1_pciexpress_cra_waitrequest),   //                   .waitrequest
		.cra_irq_irq                        (),                                               //            cra_irq.irq
		.rxm_irq_irq                        (pciexpress_rxm_irq_irq),                         //            rxm_irq.irq
		.rx_in_rx_datain_0                  (pciexpress_rx_in_rx_datain_0),                   //              rx_in.rx_datain_0
		.tx_out_tx_dataout_0                (pciexpress_tx_out_tx_dataout_0),                 //             tx_out.tx_dataout_0
		.reconfig_togxb_data                (pciexpress_reconfig_togxb_data),                 //     reconfig_togxb.data
		.reconfig_gxbclk_clk                (pll_c0_clk),                                     //    reconfig_gxbclk.clk
		.reconfig_fromgxb_0_data            (pciexpress_reconfig_fromgxb_0_data),             // reconfig_fromgxb_0.data
		.fixedclk_clk                       (pciexpress_pcie_core_clk_clk)                    //           fixedclk.clk
	);

	Architectire_PLL pll (
		.clk       (clk_clk),                            //       inclk_interface.clk
		.reset     (rst_controller_003_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                                   //             pll_slave.read
		.write     (),                                   //                      .write
		.address   (),                                   //                      .address
		.readdata  (),                                   //                      .readdata
		.writedata (),                                   //                      .writedata
		.c0        (pll_c0_clk),                         //                    c0.clk
		.c1        (clockbridge_out_clk),                //                    c1.clk
		.areset    (),                                   //        areset_conduit.export
		.locked    (),                                   //        locked_conduit.export
		.phasedone ()                                    //     phasedone_conduit.export
	);

	Architectire_Response response (
		.clk      (pciexpress_pcie_core_clk_clk),           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_response_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_response_s1_readdata), //                    .readdata
		.in_port  (response_export)                         // external_connection.export
	);

	Architectire_SGDMA sgdma (
		.clk                           (pciexpress_pcie_core_clk_clk),           //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),        //            reset.reset_n
		.csr_chipselect                (mm_interconnect_1_sgdma_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_1_sgdma_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_1_sgdma_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_1_sgdma_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_1_sgdma_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_1_sgdma_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),               //          csr_irq.irq
		.m_read_readdata               (sgdma_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_m_read_read),                      //                 .read
		.m_write_waitrequest           (sgdma_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (sgdma_m_write_address),                  //                 .address
		.m_write_write                 (sgdma_m_write_write),                    //                 .write
		.m_write_writedata             (sgdma_m_write_writedata),                //                 .writedata
		.m_write_byteenable            (sgdma_m_write_byteenable)                //                 .byteenable
	);

	Architectire_mm_interconnect_0 mm_interconnect_0 (
		.PCIExpress_pcie_core_clk_clk                                   (pciexpress_pcie_core_clk_clk),                  //                                 PCIExpress_pcie_core_clk.clk
		.PCIExpress_bar1_0_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),            // PCIExpress_bar1_0_translator_reset_reset_bridge_in_reset.reset
		.SGDMA_reset_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),                //                        SGDMA_reset_reset_bridge_in_reset.reset
		.PCIExpress_bar1_0_address                                      (pciexpress_bar1_0_address),                     //                                        PCIExpress_bar1_0.address
		.PCIExpress_bar1_0_waitrequest                                  (pciexpress_bar1_0_waitrequest),                 //                                                         .waitrequest
		.PCIExpress_bar1_0_burstcount                                   (pciexpress_bar1_0_burstcount),                  //                                                         .burstcount
		.PCIExpress_bar1_0_byteenable                                   (pciexpress_bar1_0_byteenable),                  //                                                         .byteenable
		.PCIExpress_bar1_0_read                                         (pciexpress_bar1_0_read),                        //                                                         .read
		.PCIExpress_bar1_0_readdata                                     (pciexpress_bar1_0_readdata),                    //                                                         .readdata
		.PCIExpress_bar1_0_readdatavalid                                (pciexpress_bar1_0_readdatavalid),               //                                                         .readdatavalid
		.PCIExpress_bar1_0_write                                        (pciexpress_bar1_0_write),                       //                                                         .write
		.PCIExpress_bar1_0_writedata                                    (pciexpress_bar1_0_writedata),                   //                                                         .writedata
		.SGDMA_m_write_address                                          (sgdma_m_write_address),                         //                                            SGDMA_m_write.address
		.SGDMA_m_write_waitrequest                                      (sgdma_m_write_waitrequest),                     //                                                         .waitrequest
		.SGDMA_m_write_byteenable                                       (sgdma_m_write_byteenable),                      //                                                         .byteenable
		.SGDMA_m_write_write                                            (sgdma_m_write_write),                           //                                                         .write
		.SGDMA_m_write_writedata                                        (sgdma_m_write_writedata),                       //                                                         .writedata
		.ControlSignal_s1_address                                       (mm_interconnect_0_controlsignal_s1_address),    //                                         ControlSignal_s1.address
		.ControlSignal_s1_write                                         (mm_interconnect_0_controlsignal_s1_write),      //                                                         .write
		.ControlSignal_s1_readdata                                      (mm_interconnect_0_controlsignal_s1_readdata),   //                                                         .readdata
		.ControlSignal_s1_writedata                                     (mm_interconnect_0_controlsignal_s1_writedata),  //                                                         .writedata
		.ControlSignal_s1_chipselect                                    (mm_interconnect_0_controlsignal_s1_chipselect), //                                                         .chipselect
		.FIFO_Memory_in_address                                         (mm_interconnect_0_fifo_memory_in_address),      //                                           FIFO_Memory_in.address
		.FIFO_Memory_in_write                                           (mm_interconnect_0_fifo_memory_in_write),        //                                                         .write
		.FIFO_Memory_in_writedata                                       (mm_interconnect_0_fifo_memory_in_writedata),    //                                                         .writedata
		.FIFO_Memory_in_waitrequest                                     (mm_interconnect_0_fifo_memory_in_waitrequest),  //                                                         .waitrequest
		.Response_s1_address                                            (mm_interconnect_0_response_s1_address),         //                                              Response_s1.address
		.Response_s1_readdata                                           (mm_interconnect_0_response_s1_readdata)         //                                                         .readdata
	);

	Architectire_mm_interconnect_1 mm_interconnect_1 (
		.PCIExpress_pcie_core_clk_clk                                 (pciexpress_pcie_core_clk_clk),                 //                               PCIExpress_pcie_core_clk.clk
		.PCIExpress_bar2_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),           // PCIExpress_bar2_translator_reset_reset_bridge_in_reset.reset
		.SGDMA_reset_reset_bridge_in_reset_reset                      (rst_controller_reset_out_reset),               //                      SGDMA_reset_reset_bridge_in_reset.reset
		.PCIExpress_bar2_address                                      (pciexpress_bar2_address),                      //                                        PCIExpress_bar2.address
		.PCIExpress_bar2_waitrequest                                  (pciexpress_bar2_waitrequest),                  //                                                       .waitrequest
		.PCIExpress_bar2_burstcount                                   (pciexpress_bar2_burstcount),                   //                                                       .burstcount
		.PCIExpress_bar2_byteenable                                   (pciexpress_bar2_byteenable),                   //                                                       .byteenable
		.PCIExpress_bar2_read                                         (pciexpress_bar2_read),                         //                                                       .read
		.PCIExpress_bar2_readdata                                     (pciexpress_bar2_readdata),                     //                                                       .readdata
		.PCIExpress_bar2_readdatavalid                                (pciexpress_bar2_readdatavalid),                //                                                       .readdatavalid
		.PCIExpress_bar2_write                                        (pciexpress_bar2_write),                        //                                                       .write
		.PCIExpress_bar2_writedata                                    (pciexpress_bar2_writedata),                    //                                                       .writedata
		.PCIExpress_cra_address                                       (mm_interconnect_1_pciexpress_cra_address),     //                                         PCIExpress_cra.address
		.PCIExpress_cra_write                                         (mm_interconnect_1_pciexpress_cra_write),       //                                                       .write
		.PCIExpress_cra_read                                          (mm_interconnect_1_pciexpress_cra_read),        //                                                       .read
		.PCIExpress_cra_readdata                                      (mm_interconnect_1_pciexpress_cra_readdata),    //                                                       .readdata
		.PCIExpress_cra_writedata                                     (mm_interconnect_1_pciexpress_cra_writedata),   //                                                       .writedata
		.PCIExpress_cra_byteenable                                    (mm_interconnect_1_pciexpress_cra_byteenable),  //                                                       .byteenable
		.PCIExpress_cra_waitrequest                                   (mm_interconnect_1_pciexpress_cra_waitrequest), //                                                       .waitrequest
		.PCIExpress_cra_chipselect                                    (mm_interconnect_1_pciexpress_cra_chipselect),  //                                                       .chipselect
		.SGDMA_csr_address                                            (mm_interconnect_1_sgdma_csr_address),          //                                              SGDMA_csr.address
		.SGDMA_csr_write                                              (mm_interconnect_1_sgdma_csr_write),            //                                                       .write
		.SGDMA_csr_read                                               (mm_interconnect_1_sgdma_csr_read),             //                                                       .read
		.SGDMA_csr_readdata                                           (mm_interconnect_1_sgdma_csr_readdata),         //                                                       .readdata
		.SGDMA_csr_writedata                                          (mm_interconnect_1_sgdma_csr_writedata),        //                                                       .writedata
		.SGDMA_csr_chipselect                                         (mm_interconnect_1_sgdma_csr_chipselect)        //                                                       .chipselect
	);

	Architectire_mm_interconnect_2 mm_interconnect_2 (
		.PCIExpress_pcie_core_clk_clk                                (pciexpress_pcie_core_clk_clk),                   //                              PCIExpress_pcie_core_clk.clk
		.PCIExpress_txs_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),             // PCIExpress_txs_translator_reset_reset_bridge_in_reset.reset
		.SGDMA_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),                 //                     SGDMA_reset_reset_bridge_in_reset.reset
		.SGDMA_descriptor_read_address                               (sgdma_descriptor_read_address),                  //                                 SGDMA_descriptor_read.address
		.SGDMA_descriptor_read_waitrequest                           (sgdma_descriptor_read_waitrequest),              //                                                      .waitrequest
		.SGDMA_descriptor_read_read                                  (sgdma_descriptor_read_read),                     //                                                      .read
		.SGDMA_descriptor_read_readdata                              (sgdma_descriptor_read_readdata),                 //                                                      .readdata
		.SGDMA_descriptor_read_readdatavalid                         (sgdma_descriptor_read_readdatavalid),            //                                                      .readdatavalid
		.SGDMA_descriptor_write_address                              (sgdma_descriptor_write_address),                 //                                SGDMA_descriptor_write.address
		.SGDMA_descriptor_write_waitrequest                          (sgdma_descriptor_write_waitrequest),             //                                                      .waitrequest
		.SGDMA_descriptor_write_write                                (sgdma_descriptor_write_write),                   //                                                      .write
		.SGDMA_descriptor_write_writedata                            (sgdma_descriptor_write_writedata),               //                                                      .writedata
		.SGDMA_m_read_address                                        (sgdma_m_read_address),                           //                                          SGDMA_m_read.address
		.SGDMA_m_read_waitrequest                                    (sgdma_m_read_waitrequest),                       //                                                      .waitrequest
		.SGDMA_m_read_read                                           (sgdma_m_read_read),                              //                                                      .read
		.SGDMA_m_read_readdata                                       (sgdma_m_read_readdata),                          //                                                      .readdata
		.SGDMA_m_read_readdatavalid                                  (sgdma_m_read_readdatavalid),                     //                                                      .readdatavalid
		.PCIExpress_txs_address                                      (mm_interconnect_2_pciexpress_txs_address),       //                                        PCIExpress_txs.address
		.PCIExpress_txs_write                                        (mm_interconnect_2_pciexpress_txs_write),         //                                                      .write
		.PCIExpress_txs_read                                         (mm_interconnect_2_pciexpress_txs_read),          //                                                      .read
		.PCIExpress_txs_readdata                                     (mm_interconnect_2_pciexpress_txs_readdata),      //                                                      .readdata
		.PCIExpress_txs_writedata                                    (mm_interconnect_2_pciexpress_txs_writedata),     //                                                      .writedata
		.PCIExpress_txs_burstcount                                   (mm_interconnect_2_pciexpress_txs_burstcount),    //                                                      .burstcount
		.PCIExpress_txs_byteenable                                   (mm_interconnect_2_pciexpress_txs_byteenable),    //                                                      .byteenable
		.PCIExpress_txs_readdatavalid                                (mm_interconnect_2_pciexpress_txs_readdatavalid), //                                                      .readdatavalid
		.PCIExpress_txs_waitrequest                                  (mm_interconnect_2_pciexpress_txs_waitrequest),   //                                                      .waitrequest
		.PCIExpress_txs_chipselect                                   (mm_interconnect_2_pciexpress_txs_chipselect)     //                                                      .chipselect
	);

	Architectire_irq_mapper irq_mapper (
		.clk           (pciexpress_pcie_core_clk_clk),       //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (pciexpress_rxm_irq_irq)              //    sender.irq
	);

	Architectire_avalon_st_adapter #(
		.inBitsPerSymbol (32),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (8),
		.inErrorWidth    (8),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (1),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (pciexpress_pcie_core_clk_clk),          // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (fifo_memory_out_data),                  //     in_0.data
		.in_0_valid          (fifo_memory_out_valid),                 //         .valid
		.in_0_ready          (fifo_memory_out_ready),                 //         .ready
		.in_0_startofpacket  (fifo_memory_out_startofpacket),         //         .startofpacket
		.in_0_endofpacket    (fifo_memory_out_endofpacket),           //         .endofpacket
		.in_0_error          (fifo_memory_out_error),                 //         .error
		.in_0_channel        (fifo_memory_out_channel),               //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)    //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                    // reset_in0.reset
		.reset_in1      (~pciexpress_pcie_core_reset_reset), // reset_in1.reset
		.clk            (pciexpress_pcie_core_clk_clk),      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_req      (),                                  // (terminated)
		.reset_req_in0  (1'b0),                              // (terminated)
		.reset_req_in1  (1'b0),                              // (terminated)
		.reset_in2      (1'b0),                              // (terminated)
		.reset_req_in2  (1'b0),                              // (terminated)
		.reset_in3      (1'b0),                              // (terminated)
		.reset_req_in3  (1'b0),                              // (terminated)
		.reset_in4      (1'b0),                              // (terminated)
		.reset_req_in4  (1'b0),                              // (terminated)
		.reset_in5      (1'b0),                              // (terminated)
		.reset_req_in5  (1'b0),                              // (terminated)
		.reset_in6      (1'b0),                              // (terminated)
		.reset_req_in6  (1'b0),                              // (terminated)
		.reset_in7      (1'b0),                              // (terminated)
		.reset_req_in7  (1'b0),                              // (terminated)
		.reset_in8      (1'b0),                              // (terminated)
		.reset_req_in8  (1'b0),                              // (terminated)
		.reset_in9      (1'b0),                              // (terminated)
		.reset_req_in9  (1'b0),                              // (terminated)
		.reset_in10     (1'b0),                              // (terminated)
		.reset_req_in10 (1'b0),                              // (terminated)
		.reset_in11     (1'b0),                              // (terminated)
		.reset_req_in11 (1'b0),                              // (terminated)
		.reset_in12     (1'b0),                              // (terminated)
		.reset_req_in12 (1'b0),                              // (terminated)
		.reset_in13     (1'b0),                              // (terminated)
		.reset_req_in13 (1'b0),                              // (terminated)
		.reset_in14     (1'b0),                              // (terminated)
		.reset_req_in14 (1'b0),                              // (terminated)
		.reset_in15     (1'b0),                              // (terminated)
		.reset_req_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~pciexpress_pcie_core_reset_reset),  // reset_in0.reset
		.clk            (pciexpress_pcie_core_clk_clk),       //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~pciexpress_pcie_core_reset_reset),  // reset_in1.reset
		.clk            (clockbridge_out_clk),                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
